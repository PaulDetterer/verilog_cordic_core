module tb_fdc();
//Instantiate the contoll signals
//Instantiate evaluation signals
//Generate control signals
//Instantiate dut
endmodule
